module t_Lab2_ripple_borrow_4_bit_sub;
	wire[3:0] D;
	wire B;
	reg[3:0] x,y;
	reg z;
	Lab2_ripple_borrow_4_bit_sub M1(D,B,x,y,z);
	initial begin
		x=4'b1101;y=4'b0101;z=1'b0;
	    #20	x=4'b1101;y=4'b0101;z=1'b1;
	    #20 x=4'b0101;y=4'b1101;z=1'b0;
	    #20 x=4'b0101;y=4'b1101;z=1'b1;
	    #20 x=4'b0101;y=4'b0101;z=1'b0;
	    #20	x=4'b1101;y=4'b1101;z=1'b1;
	end
	initial #200 $finish;
endmodule